
module Test;

	// Inputs
	reg [31:0] A;
	reg [31:0] B;
	reg Cin;
	reg [2:0] opcode; 
	// Outputs
	wire [31:0] Out;
	
	// Instantiate the Unit Under Test (UUT)
	FP_Adder_Sub uut (
		.A(A), 
		.B(B), 
		.Cin(Cin),
		.Out(Out),
		.opcode(opcode)
	);

	initial begin
		// Initialize Inputs
		A = 0;
		B = 0;
		Cin = 0;
		opcode = 0;
		// Wait 200 ns for global reset to finish
		#200;
       	 A=32'b01000001001101100000000000000000;//11.375
		 B=32'b01000000101100100000010000011001;//5.56300
		 Cin = 0;
		 opcode = 0;
		 //SUM=16.938
		 $monitor("Output:  %b ",Out);

		#200;
       	 A=32'b11000001001101100000000000000000;//11.375
		 B=32'b11000000101100100000010000011001;//5.56300
		 Cin = 0;
		 //SUM=16.938
		 $monitor("Output:  %b ",Out); 

	 	 #200;
       	 A=32'b01000001001101100000000000000000;//11.375
		 B=32'b11000000101100100000010000011001;//5.56300
		 Cin = 0;
		 //SUM=16.938
		 $monitor("Output:  %b ",Out);	

		 #200;
       	 A=32'b11000001001101100000000000000000;//11.375
		 B=32'b01000000101100100000010000011001;//5.56300
		 Cin = 0;
		 //SUM=16.938
		 $monitor("Output:  %b ",Out);




		#200 
		 B=32'b01000010011011111110101001111111;//59.979
		 A=32'b01000000110100000000000000000000;//6.5
		 Cin = 0;
		 opcode = 3'b001;
		 //SUM=66.479
		 $monitor("Output:  %b ",Out);
		 
		

		#200 
		 B=32'b11000010011011111110101001111111;//59.979
		 A=32'b11000000110100000000000000000000;//6.5
		 Cin = 0;
//		 opcode = 0;
		 //SUM=66.479
		 $monitor("Output:  %b ",Out);

		#200 
		 B=32'b01000010011011111110101001111111;//59.979
		 A=32'b11000000110100000000000000000000;//6.5
		 Cin = 0;
		 //SUM=66.479
		 $monitor("Output:  %b ",Out);

		#200 
		 B=32'b11000010011011111110101001111111;//59.979
		 A=32'b01000000110100000000000000000000;//6.5
		 Cin = 0;
		 //SUM=66.479
		 $monitor("Output:  %b ",Out);









		#200 
		 A=32'b01000100011110100010000000000000;//1000.5
		 B=32'b01000100011101010110100111011011;//981.654
		 Cin = 0;
		 //SUM=1982.1539
		 $monitor("Output:  %b ",Out);
		 
		 
		#200
		 A=32'b01000100000010010111111100101011;//549.987
		 B=32'b01000000101100100000010000011001;//5.563
		 Cin = 0;
		 //SUM=555.499
		 $monitor("Output:  %b ",Out);
		  
		
	end
      
endmodule
